
/***********************************************************************
  $FILENAME    : async_fifo_pkg.svh

  $TITLE       : Package definition

  $DATE        : 11 Nov 2017

  $VERSION     : 1.0.0

  $DESCRIPTION : 

Code is from: https://github.com/akzare/Async_FIFO_Verification
Verification test case for an asynchronous FIFO based on Systemverilog Object Oriented concepts and also UVM. The general architecture and implementation of the code has been taken from the UVM primer (Ray Salemi):

https://github.com/rdsalemi/uvmprimer

However the presented verification code in this test case is manipulated to be fitted for the special use case of an asynchronous FIFO.

The RTL source code for the asynchronous FIFO is taken from (Jason Yu):

http://www.verilogpro.com/asynchronous-fifo-design/

Which takes the Asynchronous FIFO design in SystemVerilog translated from Verilog to SystemVerilog, based on Cliff Cumming's Simulation and Synthesis Techniques for Asynchronous FIFO Design
http://www.sunburst-design.com/papers/CummingsSNUG2002SJ_FIFO1.pdf

************************************************************************/


package async_fifo_pkg;

  // FIFO Data Bus Width
  parameter FIFO_DATA_WIDTH = 8;
  // FIFO Address Bus Width
  parameter FIFO_MEM_ADDR_WIDTH = 4;

  `include "coverage.svh"
  `include "tester.svh"
  `include "scoreboard.svh"
  `include "tb.svh"

endpackage : async_fifo_pkg