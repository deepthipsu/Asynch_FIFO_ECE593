package definitions;

parameter [3:0] ADDRSIZE = 4'd10;
parameter [3:0] DATASIZE = 4'd8;
logic [1:0] wr_clk = 2;


endpackage
