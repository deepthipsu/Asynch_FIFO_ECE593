package definitions;

parameter [3:0] ADDRSIZE = 4'd9;
logic [1:0] wr_clk = 2;


endpackage
