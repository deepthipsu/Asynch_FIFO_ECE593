//
//
//

module Asynch_FIFO ();

endmodule
