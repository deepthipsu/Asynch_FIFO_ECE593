package definitions;

parameter ADDRSIZE = 10;
parameter DATASIZE = 8;
//parameter DEPTH = 333;
parameter WRITE_PERIOD = 2; // Number of clock cycles between successive writes
parameter READ_PERIOD = 1; // Number of clock cycles between successive reads
parameter BURST_LENGTH = 1024; // Burst length

endpackage
